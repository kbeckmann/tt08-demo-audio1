/*
 * Copyright (c) 2024 Konrad Beckmann
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_vga_example(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,   // Dedicated outputs
  input  wire [7:0] uio_in,   // IOs: Input path
  output wire [7:0] uio_out,  // IOs: Output path
  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
  input  wire       ena,      // always 1 when the design is powered, so you can ignore it
  input  wire       clk,      // clock
  input  wire       rst_n     // reset_n - low to reset
);

  // Audio signals
  wire audio_out;
  wire [15:0] audio_sample;

  // TinyVGA PMOD
  // assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};
  assign uo_out = 8'b00000000;

  // Audio PMOD
  assign uio_out = {audio_out, 7'b0000000};
  assign uio_oe = 8'b10000000;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in, uio_in};

  reg [10:0] counter;

// Audio start
  pdm #(.N(16)) pdm_gen(
    .clk(clk),
    .rst_n(rst_n),
    .pdm_in(audio_sample),
    .pdm_out(audio_out)
  );

  // ROM
  wire [8:0] rom_addr;
  reg  [8:0] rom_addr_r;
  reg  [7:0] rom_data_r;
  reg  [7:0] rom_content[512];

  initial begin
    rom_content[0] = 8'hB5;
    rom_content[1] = 8'h02;
    rom_content[2] = 8'h24;
    rom_content[3] = 8'h87;
    rom_content[4] = 8'h29;
    rom_content[5] = 8'h07;
    rom_content[6] = 8'hB5;
    rom_content[7] = 8'hC0;
    rom_content[8] = 8'hDB;
    rom_content[9] = 8'h6B;
    rom_content[10] = 8'hA6;
    rom_content[11] = 8'h59;
    rom_content[12] = 8'h37;
    rom_content[13] = 8'h8E;
    rom_content[14] = 8'hD7;
    rom_content[15] = 8'h00;
    rom_content[16] = 8'hBC;
    rom_content[17] = 8'hBC;
    rom_content[18] = 8'h58;
    rom_content[19] = 8'hDB;
    rom_content[20] = 8'hFD;
    rom_content[21] = 8'h49;
    rom_content[22] = 8'h0F;
    rom_content[23] = 8'h63;
    rom_content[24] = 8'h9B;
    rom_content[25] = 8'hA6;
    rom_content[26] = 8'h22;
    rom_content[27] = 8'hF6;
    rom_content[28] = 8'h7A;
    rom_content[29] = 8'h28;
    rom_content[30] = 8'hCB;
    rom_content[31] = 8'hE9;
    rom_content[32] = 8'h1B;
    rom_content[33] = 8'hCE;
    rom_content[34] = 8'hA8;
    rom_content[35] = 8'h37;
    rom_content[36] = 8'hA3;
    rom_content[37] = 8'hF6;
    rom_content[38] = 8'h05;
    rom_content[39] = 8'hF2;
    rom_content[40] = 8'h95;
    rom_content[41] = 8'hA8;
    rom_content[42] = 8'hBA;
    rom_content[43] = 8'h55;
    rom_content[44] = 8'h65;
    rom_content[45] = 8'hD9;
    rom_content[46] = 8'h5A;
    rom_content[47] = 8'h8B;
    rom_content[48] = 8'h09;
    rom_content[49] = 8'h72;
    rom_content[50] = 8'h57;
    rom_content[51] = 8'hCA;
    rom_content[52] = 8'h46;
    rom_content[53] = 8'hD4;
    rom_content[54] = 8'hC8;
    rom_content[55] = 8'hCB;
    rom_content[56] = 8'h7B;
    rom_content[57] = 8'h3D;
    rom_content[58] = 8'h27;
    rom_content[59] = 8'hB0;
    rom_content[60] = 8'hF1;
    rom_content[61] = 8'hFF;
    rom_content[62] = 8'hE5;
    rom_content[63] = 8'hE3;
    rom_content[64] = 8'hF6;
    rom_content[65] = 8'h1D;
    rom_content[66] = 8'h2F;
    rom_content[67] = 8'h45;
    rom_content[68] = 8'hB3;
    rom_content[69] = 8'hC2;
    rom_content[70] = 8'h06;
    rom_content[71] = 8'hCA;
    rom_content[72] = 8'hDD;
    rom_content[73] = 8'h0F;
    rom_content[74] = 8'h10;
    rom_content[75] = 8'hEA;
    rom_content[76] = 8'hB1;
    rom_content[77] = 8'h72;
    rom_content[78] = 8'hD4;
    rom_content[79] = 8'h97;
    rom_content[80] = 8'hA9;
    rom_content[81] = 8'hDC;
    rom_content[82] = 8'h3D;
    rom_content[83] = 8'h17;
    rom_content[84] = 8'h58;
    rom_content[85] = 8'hCB;
    rom_content[86] = 8'h0B;
    rom_content[87] = 8'hF7;
    rom_content[88] = 8'h2F;
    rom_content[89] = 8'hD9;
    rom_content[90] = 8'hF6;
    rom_content[91] = 8'h2F;
    rom_content[92] = 8'hD8;
    rom_content[93] = 8'h5C;
    rom_content[94] = 8'h4C;
    rom_content[95] = 8'hA9;
    rom_content[96] = 8'h1E;
    rom_content[97] = 8'h79;
    rom_content[98] = 8'hF9;
    rom_content[99] = 8'hD2;
    rom_content[100] = 8'h7E;
    rom_content[101] = 8'h0A;
    rom_content[102] = 8'hC1;
    rom_content[103] = 8'hFC;
    rom_content[104] = 8'h2F;
    rom_content[105] = 8'hD6;
    rom_content[106] = 8'hB2;
    rom_content[107] = 8'hF6;
    rom_content[108] = 8'hC9;
    rom_content[109] = 8'hDF;
    rom_content[110] = 8'h09;
    rom_content[111] = 8'h7E;
    rom_content[112] = 8'hE0;
    rom_content[113] = 8'hD9;
    rom_content[114] = 8'h43;
    rom_content[115] = 8'hB2;
    rom_content[116] = 8'h98;
    rom_content[117] = 8'hC6;
    rom_content[118] = 8'h6F;
    rom_content[119] = 8'hB9;
    rom_content[120] = 8'hEE;
    rom_content[121] = 8'h86;
    rom_content[122] = 8'hAB;
    rom_content[123] = 8'h43;
    rom_content[124] = 8'hC7;
    rom_content[125] = 8'h03;
    rom_content[126] = 8'hE1;
    rom_content[127] = 8'h3C;
    rom_content[128] = 8'h93;
    rom_content[129] = 8'hCD;
    rom_content[130] = 8'h78;
    rom_content[131] = 8'h03;
    rom_content[132] = 8'h79;
    rom_content[133] = 8'h71;
    rom_content[134] = 8'hAA;
    rom_content[135] = 8'hC5;
    rom_content[136] = 8'hF2;
    rom_content[137] = 8'h6E;
    rom_content[138] = 8'hFD;
    rom_content[139] = 8'hFC;
    rom_content[140] = 8'hA9;
    rom_content[141] = 8'h82;
    rom_content[142] = 8'h91;
    rom_content[143] = 8'h74;
    rom_content[144] = 8'h46;
    rom_content[145] = 8'h1E;
    rom_content[146] = 8'hD5;
    rom_content[147] = 8'h2E;
    rom_content[148] = 8'h40;
    rom_content[149] = 8'h4B;
    rom_content[150] = 8'h43;
    rom_content[151] = 8'h6C;
    rom_content[152] = 8'h8A;
    rom_content[153] = 8'hE2;
    rom_content[154] = 8'h93;
    rom_content[155] = 8'hA8;
    rom_content[156] = 8'h53;
    rom_content[157] = 8'h69;
    rom_content[158] = 8'hB1;
    rom_content[159] = 8'hC1;
    rom_content[160] = 8'h76;
    rom_content[161] = 8'h7A;
    rom_content[162] = 8'hA0;
    rom_content[163] = 8'h36;
    rom_content[164] = 8'h39;
    rom_content[165] = 8'h15;
    rom_content[166] = 8'hF6;
    rom_content[167] = 8'hCB;
    rom_content[168] = 8'h84;
    rom_content[169] = 8'hFF;
    rom_content[170] = 8'h3E;
    rom_content[171] = 8'h14;
    rom_content[172] = 8'hEC;
    rom_content[173] = 8'h18;
    rom_content[174] = 8'hBB;
    rom_content[175] = 8'h18;
    rom_content[176] = 8'hCD;
    rom_content[177] = 8'h0B;
    rom_content[178] = 8'h30;
    rom_content[179] = 8'hE1;
    rom_content[180] = 8'h83;
    rom_content[181] = 8'hE9;
    rom_content[182] = 8'h2C;
    rom_content[183] = 8'hAD;
    rom_content[184] = 8'h69;
    rom_content[185] = 8'hD0;
    rom_content[186] = 8'hEB;
    rom_content[187] = 8'h9B;
    rom_content[188] = 8'hF9;
    rom_content[189] = 8'hBD;
    rom_content[190] = 8'hD0;
    rom_content[191] = 8'hDC;
    rom_content[192] = 8'h5C;
    rom_content[193] = 8'h1E;
    rom_content[194] = 8'h11;
    rom_content[195] = 8'h34;
    rom_content[196] = 8'h98;
    rom_content[197] = 8'h95;
    rom_content[198] = 8'h8E;
    rom_content[199] = 8'hA3;
    rom_content[200] = 8'hD5;
    rom_content[201] = 8'h0D;
    rom_content[202] = 8'h67;
    rom_content[203] = 8'hD0;
    rom_content[204] = 8'hE9;
    rom_content[205] = 8'hAF;
    rom_content[206] = 8'hDA;
    rom_content[207] = 8'h79;
    rom_content[208] = 8'hE8;
    rom_content[209] = 8'h6B;
    rom_content[210] = 8'h0A;
    rom_content[211] = 8'h9E;
    rom_content[212] = 8'h3B;
    rom_content[213] = 8'h63;
    rom_content[214] = 8'hFD;
    rom_content[215] = 8'h0A;
    rom_content[216] = 8'hB1;
    rom_content[217] = 8'h9A;
    rom_content[218] = 8'hA9;
    rom_content[219] = 8'h93;
    rom_content[220] = 8'h77;
    rom_content[221] = 8'h4A;
    rom_content[222] = 8'h16;
    rom_content[223] = 8'h94;
    rom_content[224] = 8'h43;
    rom_content[225] = 8'h3E;
    rom_content[226] = 8'hF2;
    rom_content[227] = 8'hAF;
    rom_content[228] = 8'h1B;
    rom_content[229] = 8'h16;
    rom_content[230] = 8'h16;
    rom_content[231] = 8'hBD;
    rom_content[232] = 8'h71;
    rom_content[233] = 8'h85;
    rom_content[234] = 8'h6D;
    rom_content[235] = 8'h88;
    rom_content[236] = 8'h09;
    rom_content[237] = 8'h4C;
    rom_content[238] = 8'h6D;
    rom_content[239] = 8'h3F;
    rom_content[240] = 8'hA5;
    rom_content[241] = 8'hC9;
    rom_content[242] = 8'hA3;
    rom_content[243] = 8'h0A;
    rom_content[244] = 8'h96;
    rom_content[245] = 8'h52;
    rom_content[246] = 8'h8C;
    rom_content[247] = 8'h7B;
    rom_content[248] = 8'hFA;
    rom_content[249] = 8'h80;
    rom_content[250] = 8'hDD;
    rom_content[251] = 8'hB3;
    rom_content[252] = 8'h77;
    rom_content[253] = 8'h2C;
    rom_content[254] = 8'hC4;
    rom_content[255] = 8'hE6;
    rom_content[256] = 8'hB5;
    rom_content[257] = 8'h3B;
    rom_content[258] = 8'hE6;
    rom_content[259] = 8'hB1;
    rom_content[260] = 8'hDB;
    rom_content[261] = 8'h77;
    rom_content[262] = 8'h42;
    rom_content[263] = 8'h7E;
    rom_content[264] = 8'h1C;
    rom_content[265] = 8'hAC;
    rom_content[266] = 8'hEB;
    rom_content[267] = 8'hEF;
    rom_content[268] = 8'h61;
    rom_content[269] = 8'hD6;
    rom_content[270] = 8'hE2;
    rom_content[271] = 8'hF6;
    rom_content[272] = 8'h08;
    rom_content[273] = 8'h40;
    rom_content[274] = 8'h9F;
    rom_content[275] = 8'h04;
    rom_content[276] = 8'h52;
    rom_content[277] = 8'h23;
    rom_content[278] = 8'h90;
    rom_content[279] = 8'hDF;
    rom_content[280] = 8'h49;
    rom_content[281] = 8'hBF;
    rom_content[282] = 8'h55;
    rom_content[283] = 8'hE9;
    rom_content[284] = 8'h4E;
    rom_content[285] = 8'h99;
    rom_content[286] = 8'h67;
    rom_content[287] = 8'hE4;
    rom_content[288] = 8'hFD;
    rom_content[289] = 8'h35;
    rom_content[290] = 8'h34;
    rom_content[291] = 8'h8C;
    rom_content[292] = 8'h51;
    rom_content[293] = 8'h0A;
    rom_content[294] = 8'h5C;
    rom_content[295] = 8'h46;
    rom_content[296] = 8'hE3;
    rom_content[297] = 8'h19;
    rom_content[298] = 8'hB8;
    rom_content[299] = 8'h41;
    rom_content[300] = 8'h42;
    rom_content[301] = 8'h35;
    rom_content[302] = 8'hA3;
    rom_content[303] = 8'h01;
    rom_content[304] = 8'h5C;
    rom_content[305] = 8'h86;
    rom_content[306] = 8'h8A;
    rom_content[307] = 8'hD2;
    rom_content[308] = 8'h87;
    rom_content[309] = 8'hFF;
    rom_content[310] = 8'h20;
    rom_content[311] = 8'hA6;
    rom_content[312] = 8'hEC;
    rom_content[313] = 8'hF8;
    rom_content[314] = 8'hF2;
    rom_content[315] = 8'hA8;
    rom_content[316] = 8'h2E;
    rom_content[317] = 8'h81;
    rom_content[318] = 8'h64;
    rom_content[319] = 8'h29;
    rom_content[320] = 8'hF6;
    rom_content[321] = 8'hBC;
    rom_content[322] = 8'h11;
    rom_content[323] = 8'h5B;
    rom_content[324] = 8'hD6;
    rom_content[325] = 8'hED;
    rom_content[326] = 8'h2D;
    rom_content[327] = 8'h9E;
    rom_content[328] = 8'hFF;
    rom_content[329] = 8'h8B;
    rom_content[330] = 8'h2E;
    rom_content[331] = 8'hC7;
    rom_content[332] = 8'h42;
    rom_content[333] = 8'h9A;
    rom_content[334] = 8'h86;
    rom_content[335] = 8'h62;
    rom_content[336] = 8'h25;
    rom_content[337] = 8'h94;
    rom_content[338] = 8'h34;
    rom_content[339] = 8'h19;
    rom_content[340] = 8'hE9;
    rom_content[341] = 8'hD4;
    rom_content[342] = 8'hC7;
    rom_content[343] = 8'hA9;
    rom_content[344] = 8'hB4;
    rom_content[345] = 8'h6D;
    rom_content[346] = 8'h83;
    rom_content[347] = 8'h98;
    rom_content[348] = 8'hA8;
    rom_content[349] = 8'hC4;
    rom_content[350] = 8'h3A;
    rom_content[351] = 8'h27;
    rom_content[352] = 8'hB5;
    rom_content[353] = 8'h2A;
    rom_content[354] = 8'hEC;
    rom_content[355] = 8'h76;
    rom_content[356] = 8'h1B;
    rom_content[357] = 8'h13;
    rom_content[358] = 8'hDB;
    rom_content[359] = 8'h76;
    rom_content[360] = 8'hF7;
    rom_content[361] = 8'h4D;
    rom_content[362] = 8'hA7;
    rom_content[363] = 8'h5A;
    rom_content[364] = 8'hFB;
    rom_content[365] = 8'hB5;
    rom_content[366] = 8'h92;
    rom_content[367] = 8'h5A;
    rom_content[368] = 8'hD3;
    rom_content[369] = 8'h6D;
    rom_content[370] = 8'h18;
    rom_content[371] = 8'hA6;
    rom_content[372] = 8'h11;
    rom_content[373] = 8'hB4;
    rom_content[374] = 8'h90;
    rom_content[375] = 8'h6D;
    rom_content[376] = 8'h67;
    rom_content[377] = 8'h90;
    rom_content[378] = 8'hEE;
    rom_content[379] = 8'h89;
    rom_content[380] = 8'hB6;
    rom_content[381] = 8'hA0;
    rom_content[382] = 8'h7C;
    rom_content[383] = 8'h23;
    rom_content[384] = 8'h8F;
    rom_content[385] = 8'h4E;
    rom_content[386] = 8'hEC;
    rom_content[387] = 8'h2A;
    rom_content[388] = 8'hDC;
    rom_content[389] = 8'h15;
    rom_content[390] = 8'h5E;
    rom_content[391] = 8'h37;
    rom_content[392] = 8'h83;
    rom_content[393] = 8'h02;
    rom_content[394] = 8'h0F;
    rom_content[395] = 8'hAB;
    rom_content[396] = 8'h12;
    rom_content[397] = 8'hF9;
    rom_content[398] = 8'hAA;
    rom_content[399] = 8'h44;
    rom_content[400] = 8'h39;
    rom_content[401] = 8'hDB;
    rom_content[402] = 8'h23;
    rom_content[403] = 8'h3F;
    rom_content[404] = 8'hB3;
    rom_content[405] = 8'hB3;
    rom_content[406] = 8'h23;
    rom_content[407] = 8'hCF;
    rom_content[408] = 8'h31;
    rom_content[409] = 8'h3E;
    rom_content[410] = 8'h02;
    rom_content[411] = 8'hC6;
    rom_content[412] = 8'hD3;
    rom_content[413] = 8'h20;
    rom_content[414] = 8'h7F;
    rom_content[415] = 8'hD5;
    rom_content[416] = 8'hE9;
    rom_content[417] = 8'h76;
    rom_content[418] = 8'hA9;
    rom_content[419] = 8'h04;
    rom_content[420] = 8'h97;
    rom_content[421] = 8'hEA;
    rom_content[422] = 8'hBB;
    rom_content[423] = 8'h2E;
    rom_content[424] = 8'hE7;
    rom_content[425] = 8'hFC;
    rom_content[426] = 8'h3A;
    rom_content[427] = 8'h6E;
    rom_content[428] = 8'h0F;
    rom_content[429] = 8'hBE;
    rom_content[430] = 8'h17;
    rom_content[431] = 8'h1A;
    rom_content[432] = 8'h1C;
    rom_content[433] = 8'hE6;
    rom_content[434] = 8'hA9;
    rom_content[435] = 8'hBE;
    rom_content[436] = 8'hDB;
    rom_content[437] = 8'h82;
    rom_content[438] = 8'h4E;
    rom_content[439] = 8'h54;
    rom_content[440] = 8'hBB;
    rom_content[441] = 8'h6B;
    rom_content[442] = 8'h80;
    rom_content[443] = 8'hEB;
    rom_content[444] = 8'hF1;
    rom_content[445] = 8'hA7;
    rom_content[446] = 8'hD2;
    rom_content[447] = 8'hB1;
    rom_content[448] = 8'hB3;
    rom_content[449] = 8'h69;
    rom_content[450] = 8'h10;
    rom_content[451] = 8'h40;
    rom_content[452] = 8'h51;
    rom_content[453] = 8'h23;
    rom_content[454] = 8'h0F;
    rom_content[455] = 8'hA4;
    rom_content[456] = 8'h27;
    rom_content[457] = 8'hDA;
    rom_content[458] = 8'h4B;
    rom_content[459] = 8'h9E;
    rom_content[460] = 8'hF1;
    rom_content[461] = 8'h45;
    rom_content[462] = 8'h1E;
    rom_content[463] = 8'h9D;
    rom_content[464] = 8'h4A;
    rom_content[465] = 8'h7D;
    rom_content[466] = 8'h4B;
    rom_content[467] = 8'h40;
    rom_content[468] = 8'h7B;
    rom_content[469] = 8'h85;
    rom_content[470] = 8'h32;
    rom_content[471] = 8'h8A;
    rom_content[472] = 8'h20;
    rom_content[473] = 8'h1C;
    rom_content[474] = 8'hD4;
    rom_content[475] = 8'h66;
    rom_content[476] = 8'h15;
    rom_content[477] = 8'hEF;
    rom_content[478] = 8'hAD;
    rom_content[479] = 8'h60;
    rom_content[480] = 8'h1F;
    rom_content[481] = 8'h9E;
    rom_content[482] = 8'h2D;
    rom_content[483] = 8'hE2;
    rom_content[484] = 8'h14;
    rom_content[485] = 8'h09;
    rom_content[486] = 8'h47;
    rom_content[487] = 8'hB5;
    rom_content[488] = 8'hBD;
    rom_content[489] = 8'h65;
    rom_content[490] = 8'h8A;
    rom_content[491] = 8'hF1;
    rom_content[492] = 8'h4D;
    rom_content[493] = 8'h2F;
    rom_content[494] = 8'h34;
    rom_content[495] = 8'hE7;
    rom_content[496] = 8'h96;
    rom_content[497] = 8'hE8;
    rom_content[498] = 8'hD0;
    rom_content[499] = 8'h9C;
    rom_content[500] = 8'hCA;
    rom_content[501] = 8'hFB;
    rom_content[502] = 8'h65;
    rom_content[503] = 8'hF2;
    rom_content[504] = 8'h58;
    rom_content[505] = 8'h6E;
    rom_content[506] = 8'hFF;
    rom_content[507] = 8'h19;
    rom_content[508] = 8'h2F;
    rom_content[509] = 8'h89;
    rom_content[510] = 8'h7F;
    rom_content[511] = 8'h1D;
  end

  always @(posedge clk) begin
    if (~rst_n) begin
      rom_addr_r <= 0;
      rom_data_r <= 0;
    end else begin
      rom_addr_r <= rom_addr;
      rom_data_r <= rom_content[rom_addr_r];
    end
  end

  assign rom_addr = counter[10:2];
  assign audio_sample = {8'h00, rom_data_r};

// Audio end

  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      counter <= counter + 1;
    end
  end
  
endmodule
