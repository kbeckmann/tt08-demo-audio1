/*
 * Copyright (c) 2024 Konrad Beckmann
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_vga_example(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,   // Dedicated outputs
  input  wire [7:0] uio_in,   // IOs: Input path
  output wire [7:0] uio_out,  // IOs: Output path
  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
  input  wire       ena,      // always 1 when the design is powered, so you can ignore it
  input  wire       clk,      // clock
  input  wire       rst_n     // reset_n - low to reset
);

  // Audio signals
  wire audio_out;
  wire [15:0] audio_sample;

  // TinyVGA PMOD
  // assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};
  assign uo_out = 8'b00000000;

  // Audio PMOD
  assign uio_out = {audio_out, 7'b0000000};
  assign uio_oe = 8'b10000000;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in, uio_in};

  reg [10:0] counter;

// Audio start
  pdm #(.N(16)) pdm_gen(
    .clk(clk),
    .rst_n(rst_n),
    .pdm_in(audio_sample),
    .pdm_out(audio_out)
  );

  // ROM
  wire [8:0] rom_addr;
  reg  [8:0] rom_addr_r;
  reg  [7:0] rom_data;
  reg  [7:0] rom_data_r;

  always @(*) begin
    case (rom_addr_r)
      9'h000: rom_data = 8'h22;
      9'h001: rom_data = 8'h89;
      9'h002: rom_data = 8'h91;
      9'h003: rom_data = 8'h27;
      9'h004: rom_data = 8'h79;
      9'h005: rom_data = 8'hD2;
      9'h006: rom_data = 8'h62;
      9'h007: rom_data = 8'hAE;
      9'h008: rom_data = 8'h9F;
      9'h009: rom_data = 8'h59;
      9'h00A: rom_data = 8'h1B;
      9'h00B: rom_data = 8'h6A;
      9'h00C: rom_data = 8'hAD;
      9'h00D: rom_data = 8'h4E;
      9'h00E: rom_data = 8'hFD;
      9'h00F: rom_data = 8'h56;
      9'h010: rom_data = 8'h6A;
      9'h011: rom_data = 8'h17;
      9'h012: rom_data = 8'hE1;
      9'h013: rom_data = 8'h6E;
      9'h014: rom_data = 8'h5B;
      9'h015: rom_data = 8'h0D;
      9'h016: rom_data = 8'hFE;
      9'h017: rom_data = 8'hF6;
      9'h018: rom_data = 8'h18;
      9'h019: rom_data = 8'h60;
      9'h01A: rom_data = 8'h3A;
      9'h01B: rom_data = 8'h70;
      9'h01C: rom_data = 8'h0A;
      9'h01D: rom_data = 8'h13;
      9'h01E: rom_data = 8'hEA;
      9'h01F: rom_data = 8'hB9;
      9'h020: rom_data = 8'h36;
      9'h021: rom_data = 8'hCA;
      9'h022: rom_data = 8'hBC;
      9'h023: rom_data = 8'h8E;
      9'h024: rom_data = 8'h4A;
      9'h025: rom_data = 8'h63;
      9'h026: rom_data = 8'h59;
      9'h027: rom_data = 8'h85;
      9'h028: rom_data = 8'hE2;
      9'h029: rom_data = 8'h13;
      9'h02A: rom_data = 8'hFC;
      9'h02B: rom_data = 8'hF2;
      9'h02C: rom_data = 8'h5D;
      9'h02D: rom_data = 8'hB3;
      9'h02E: rom_data = 8'hCA;
      9'h02F: rom_data = 8'h52;
      9'h030: rom_data = 8'h2D;
      9'h031: rom_data = 8'hF2;
      9'h032: rom_data = 8'hFF;
      9'h033: rom_data = 8'h5E;
      9'h034: rom_data = 8'hA4;
      9'h035: rom_data = 8'hBD;
      9'h036: rom_data = 8'h37;
      9'h037: rom_data = 8'hDF;
      9'h038: rom_data = 8'hF0;
      9'h039: rom_data = 8'h21;
      9'h03A: rom_data = 8'h3A;
      9'h03B: rom_data = 8'h5F;
      9'h03C: rom_data = 8'hF3;
      9'h03D: rom_data = 8'hDD;
      9'h03E: rom_data = 8'h23;
      9'h03F: rom_data = 8'h20;
      9'h040: rom_data = 8'h15;
      9'h041: rom_data = 8'hCF;
      9'h042: rom_data = 8'h31;
      9'h043: rom_data = 8'hD5;
      9'h044: rom_data = 8'hE8;
      9'h045: rom_data = 8'hBD;
      9'h046: rom_data = 8'h6B;
      9'h047: rom_data = 8'h59;
      9'h048: rom_data = 8'h14;
      9'h049: rom_data = 8'h84;
      9'h04A: rom_data = 8'h12;
      9'h04B: rom_data = 8'h13;
      9'h04C: rom_data = 8'h96;
      9'h04D: rom_data = 8'hA2;
      9'h04E: rom_data = 8'h98;
      9'h04F: rom_data = 8'h60;
      9'h050: rom_data = 8'hF2;
      9'h051: rom_data = 8'h9E;
      9'h052: rom_data = 8'h78;
      9'h053: rom_data = 8'hF7;
      9'h054: rom_data = 8'h46;
      9'h055: rom_data = 8'h4D;
      9'h056: rom_data = 8'h65;
      9'h057: rom_data = 8'h06;
      9'h058: rom_data = 8'hA9;
      9'h059: rom_data = 8'h90;
      9'h05A: rom_data = 8'h49;
      9'h05B: rom_data = 8'h4B;
      9'h05C: rom_data = 8'h63;
      9'h05D: rom_data = 8'hD7;
      9'h05E: rom_data = 8'h31;
      9'h05F: rom_data = 8'hC6;
      9'h060: rom_data = 8'h4A;
      9'h061: rom_data = 8'h26;
      9'h062: rom_data = 8'h27;
      9'h063: rom_data = 8'h03;
      9'h064: rom_data = 8'h63;
      9'h065: rom_data = 8'h6B;
      9'h066: rom_data = 8'h97;
      9'h067: rom_data = 8'h47;
      9'h068: rom_data = 8'hC5;
      9'h069: rom_data = 8'h78;
      9'h06A: rom_data = 8'hCD;
      9'h06B: rom_data = 8'h20;
      9'h06C: rom_data = 8'h1F;
      9'h06D: rom_data = 8'h0A;
      9'h06E: rom_data = 8'hF0;
      9'h06F: rom_data = 8'h25;
      9'h070: rom_data = 8'h40;
      9'h071: rom_data = 8'h4D;
      9'h072: rom_data = 8'hB5;
      9'h073: rom_data = 8'h53;
      9'h074: rom_data = 8'h5C;
      9'h075: rom_data = 8'hBE;
      9'h076: rom_data = 8'h83;
      9'h077: rom_data = 8'h7B;
      9'h078: rom_data = 8'h98;
      9'h079: rom_data = 8'h03;
      9'h07A: rom_data = 8'hC5;
      9'h07B: rom_data = 8'h05;
      9'h07C: rom_data = 8'h8F;
      9'h07D: rom_data = 8'hB9;
      9'h07E: rom_data = 8'h8E;
      9'h07F: rom_data = 8'hAF;
      9'h080: rom_data = 8'hF4;
      9'h081: rom_data = 8'h06;
      9'h082: rom_data = 8'h24;
      9'h083: rom_data = 8'h86;
      9'h084: rom_data = 8'h0A;
      9'h085: rom_data = 8'h8A;
      9'h086: rom_data = 8'hF2;
      9'h087: rom_data = 8'h9C;
      9'h088: rom_data = 8'hDE;
      9'h089: rom_data = 8'h64;
      9'h08A: rom_data = 8'h92;
      9'h08B: rom_data = 8'h83;
      9'h08C: rom_data = 8'hA8;
      9'h08D: rom_data = 8'h73;
      9'h08E: rom_data = 8'h99;
      9'h08F: rom_data = 8'hFF;
      9'h090: rom_data = 8'h3E;
      9'h091: rom_data = 8'hD6;
      9'h092: rom_data = 8'hCB;
      9'h093: rom_data = 8'hF8;
      9'h094: rom_data = 8'hEB;
      9'h095: rom_data = 8'h1B;
      9'h096: rom_data = 8'hFD;
      9'h097: rom_data = 8'h28;
      9'h098: rom_data = 8'hD8;
      9'h099: rom_data = 8'hB7;
      9'h09A: rom_data = 8'h24;
      9'h09B: rom_data = 8'h06;
      9'h09C: rom_data = 8'h40;
      9'h09D: rom_data = 8'h5F;
      9'h09E: rom_data = 8'h80;
      9'h09F: rom_data = 8'h5C;
      9'h0A0: rom_data = 8'hCC;
      9'h0A1: rom_data = 8'hC8;
      9'h0A2: rom_data = 8'h0C;
      9'h0A3: rom_data = 8'h31;
      9'h0A4: rom_data = 8'hDD;
      9'h0A5: rom_data = 8'h00;
      9'h0A6: rom_data = 8'h4C;
      9'h0A7: rom_data = 8'hBA;
      9'h0A8: rom_data = 8'h03;
      9'h0A9: rom_data = 8'hC3;
      9'h0AA: rom_data = 8'hE4;
      9'h0AB: rom_data = 8'h2B;
      9'h0AC: rom_data = 8'h8E;
      9'h0AD: rom_data = 8'hBC;
      9'h0AE: rom_data = 8'h4D;
      9'h0AF: rom_data = 8'h31;
      9'h0B0: rom_data = 8'h39;
      9'h0B1: rom_data = 8'h8F;
      9'h0B2: rom_data = 8'h79;
      9'h0B3: rom_data = 8'h5C;
      9'h0B4: rom_data = 8'h85;
      9'h0B5: rom_data = 8'hEA;
      9'h0B6: rom_data = 8'h2A;
      9'h0B7: rom_data = 8'h39;
      9'h0B8: rom_data = 8'h32;
      9'h0B9: rom_data = 8'hE9;
      9'h0BA: rom_data = 8'h65;
      9'h0BB: rom_data = 8'h93;
      9'h0BC: rom_data = 8'hF2;
      9'h0BD: rom_data = 8'hB6;
      9'h0BE: rom_data = 8'h15;
      9'h0BF: rom_data = 8'h98;
      9'h0C0: rom_data = 8'hA8;
      9'h0C1: rom_data = 8'h47;
      9'h0C2: rom_data = 8'hB0;
      9'h0C3: rom_data = 8'h58;
      9'h0C4: rom_data = 8'hB5;
      9'h0C5: rom_data = 8'hFD;
      9'h0C6: rom_data = 8'hD8;
      9'h0C7: rom_data = 8'hA2;
      9'h0C8: rom_data = 8'hCC;
      9'h0C9: rom_data = 8'h14;
      9'h0CA: rom_data = 8'h7D;
      9'h0CB: rom_data = 8'h8C;
      9'h0CC: rom_data = 8'h06;
      9'h0CD: rom_data = 8'hE5;
      9'h0CE: rom_data = 8'hDA;
      9'h0CF: rom_data = 8'h21;
      9'h0D0: rom_data = 8'h4B;
      9'h0D1: rom_data = 8'h46;
      9'h0D2: rom_data = 8'h5E;
      9'h0D3: rom_data = 8'hA7;
      9'h0D4: rom_data = 8'h67;
      9'h0D5: rom_data = 8'h99;
      9'h0D6: rom_data = 8'h08;
      9'h0D7: rom_data = 8'hFB;
      9'h0D8: rom_data = 8'h06;
      9'h0D9: rom_data = 8'h05;
      9'h0DA: rom_data = 8'hF4;
      9'h0DB: rom_data = 8'h4E;
      9'h0DC: rom_data = 8'hEA;
      9'h0DD: rom_data = 8'hDE;
      9'h0DE: rom_data = 8'h77;
      9'h0DF: rom_data = 8'h29;
      9'h0E0: rom_data = 8'h71;
      9'h0E1: rom_data = 8'hE1;
      9'h0E2: rom_data = 8'h4A;
      9'h0E3: rom_data = 8'h3B;
      9'h0E4: rom_data = 8'hB9;
      9'h0E5: rom_data = 8'h2A;
      9'h0E6: rom_data = 8'hD6;
      9'h0E7: rom_data = 8'hC7;
      9'h0E8: rom_data = 8'hB3;
      9'h0E9: rom_data = 8'h94;
      9'h0EA: rom_data = 8'h23;
      9'h0EB: rom_data = 8'h56;
      9'h0EC: rom_data = 8'h67;
      9'h0ED: rom_data = 8'h4E;
      9'h0EE: rom_data = 8'hA4;
      9'h0EF: rom_data = 8'hB4;
      9'h0F0: rom_data = 8'h1C;
      9'h0F1: rom_data = 8'h80;
      9'h0F2: rom_data = 8'h3B;
      9'h0F3: rom_data = 8'hB8;
      9'h0F4: rom_data = 8'h16;
      9'h0F5: rom_data = 8'hAF;
      9'h0F6: rom_data = 8'hC9;
      9'h0F7: rom_data = 8'h29;
      9'h0F8: rom_data = 8'hFF;
      9'h0F9: rom_data = 8'h28;
      9'h0FA: rom_data = 8'hC3;
      9'h0FB: rom_data = 8'h51;
      9'h0FC: rom_data = 8'h62;
      9'h0FD: rom_data = 8'h86;
      9'h0FE: rom_data = 8'hAF;
      9'h0FF: rom_data = 8'h35;
      9'h100: rom_data = 8'h61;
      9'h101: rom_data = 8'h23;
      9'h102: rom_data = 8'h63;
      9'h103: rom_data = 8'hDE;
      9'h104: rom_data = 8'h3E;
      9'h105: rom_data = 8'hFB;
      9'h106: rom_data = 8'h75;
      9'h107: rom_data = 8'h68;
      9'h108: rom_data = 8'hD1;
      9'h109: rom_data = 8'h61;
      9'h10A: rom_data = 8'hF4;
      9'h10B: rom_data = 8'hEF;
      9'h10C: rom_data = 8'hE4;
      9'h10D: rom_data = 8'h0C;
      9'h10E: rom_data = 8'hEB;
      9'h10F: rom_data = 8'hB3;
      9'h110: rom_data = 8'hF1;
      9'h111: rom_data = 8'h80;
      9'h112: rom_data = 8'h61;
      9'h113: rom_data = 8'hA5;
      9'h114: rom_data = 8'hC1;
      9'h115: rom_data = 8'h54;
      9'h116: rom_data = 8'hF4;
      9'h117: rom_data = 8'hC6;
      9'h118: rom_data = 8'h1D;
      9'h119: rom_data = 8'hBC;
      9'h11A: rom_data = 8'hA1;
      9'h11B: rom_data = 8'h6F;
      9'h11C: rom_data = 8'h85;
      9'h11D: rom_data = 8'hEB;
      9'h11E: rom_data = 8'hE9;
      9'h11F: rom_data = 8'h5A;
      9'h120: rom_data = 8'hA2;
      9'h121: rom_data = 8'h78;
      9'h122: rom_data = 8'h02;
      9'h123: rom_data = 8'hF7;
      9'h124: rom_data = 8'h7E;
      9'h125: rom_data = 8'hAA;
      9'h126: rom_data = 8'h48;
      9'h127: rom_data = 8'hB7;
      9'h128: rom_data = 8'h17;
      9'h129: rom_data = 8'h5D;
      9'h12A: rom_data = 8'hB5;
      9'h12B: rom_data = 8'h7B;
      9'h12C: rom_data = 8'hA4;
      9'h12D: rom_data = 8'h4E;
      9'h12E: rom_data = 8'h18;
      9'h12F: rom_data = 8'hC4;
      9'h130: rom_data = 8'h92;
      9'h131: rom_data = 8'hD9;
      9'h132: rom_data = 8'hC3;
      9'h133: rom_data = 8'h09;
      9'h134: rom_data = 8'h34;
      9'h135: rom_data = 8'h7B;
      9'h136: rom_data = 8'hAB;
      9'h137: rom_data = 8'h95;
      9'h138: rom_data = 8'h82;
      9'h139: rom_data = 8'h2F;
      9'h13A: rom_data = 8'h57;
      9'h13B: rom_data = 8'h5E;
      9'h13C: rom_data = 8'hCC;
      9'h13D: rom_data = 8'hB3;
      9'h13E: rom_data = 8'hAD;
      9'h13F: rom_data = 8'h54;
      9'h140: rom_data = 8'hEB;
      9'h141: rom_data = 8'hC4;
      9'h142: rom_data = 8'h83;
      9'h143: rom_data = 8'h27;
      9'h144: rom_data = 8'hD1;
      9'h145: rom_data = 8'hA0;
      9'h146: rom_data = 8'hD5;
      9'h147: rom_data = 8'h17;
      9'h148: rom_data = 8'h0F;
      9'h149: rom_data = 8'h9F;
      9'h14A: rom_data = 8'h59;
      9'h14B: rom_data = 8'hE3;
      9'h14C: rom_data = 8'h3E;
      9'h14D: rom_data = 8'hD0;
      9'h14E: rom_data = 8'hD8;
      9'h14F: rom_data = 8'hAD;
      9'h150: rom_data = 8'h5F;
      9'h151: rom_data = 8'hD7;
      9'h152: rom_data = 8'h1C;
      9'h153: rom_data = 8'hEC;
      9'h154: rom_data = 8'hF1;
      9'h155: rom_data = 8'hEF;
      9'h156: rom_data = 8'h33;
      9'h157: rom_data = 8'hF9;
      9'h158: rom_data = 8'h46;
      9'h159: rom_data = 8'h5B;
      9'h15A: rom_data = 8'h40;
      9'h15B: rom_data = 8'h67;
      9'h15C: rom_data = 8'hDE;
      9'h15D: rom_data = 8'h4B;
      9'h15E: rom_data = 8'h51;
      9'h15F: rom_data = 8'h70;
      9'h160: rom_data = 8'h80;
      9'h161: rom_data = 8'hC7;
      9'h162: rom_data = 8'hE0;
      9'h163: rom_data = 8'h32;
      9'h164: rom_data = 8'hBB;
      9'h165: rom_data = 8'hE8;
      9'h166: rom_data = 8'h83;
      9'h167: rom_data = 8'hC2;
      9'h168: rom_data = 8'h05;
      9'h169: rom_data = 8'h9D;
      9'h16A: rom_data = 8'h89;
      9'h16B: rom_data = 8'hD4;
      9'h16C: rom_data = 8'h16;
      9'h16D: rom_data = 8'h60;
      9'h16E: rom_data = 8'hB4;
      9'h16F: rom_data = 8'h82;
      9'h170: rom_data = 8'h5F;
      9'h171: rom_data = 8'hEA;
      9'h172: rom_data = 8'h3E;
      9'h173: rom_data = 8'h3D;
      9'h174: rom_data = 8'h6A;
      9'h175: rom_data = 8'h16;
      9'h176: rom_data = 8'h24;
      9'h177: rom_data = 8'hB8;
      9'h178: rom_data = 8'h6F;
      9'h179: rom_data = 8'h20;
      9'h17A: rom_data = 8'h51;
      9'h17B: rom_data = 8'h4D;
      9'h17C: rom_data = 8'h8B;
      9'h17D: rom_data = 8'h92;
      9'h17E: rom_data = 8'hD7;
      9'h17F: rom_data = 8'h09;
      9'h180: rom_data = 8'h39;
      9'h181: rom_data = 8'h02;
      9'h182: rom_data = 8'hDD;
      9'h183: rom_data = 8'h61;
      9'h184: rom_data = 8'hFB;
      9'h185: rom_data = 8'h1C;
      9'h186: rom_data = 8'h98;
      9'h187: rom_data = 8'hD4;
      9'h188: rom_data = 8'hA4;
      9'h189: rom_data = 8'h27;
      9'h18A: rom_data = 8'hE6;
      9'h18B: rom_data = 8'h78;
      9'h18C: rom_data = 8'h88;
      9'h18D: rom_data = 8'hED;
      9'h18E: rom_data = 8'h95;
      9'h18F: rom_data = 8'h27;
      9'h190: rom_data = 8'h30;
      9'h191: rom_data = 8'h1B;
      9'h192: rom_data = 8'hBB;
      9'h193: rom_data = 8'hB2;
      9'h194: rom_data = 8'h3F;
      9'h195: rom_data = 8'h32;
      9'h196: rom_data = 8'hA7;
      9'h197: rom_data = 8'hF2;
      9'h198: rom_data = 8'hC2;
      9'h199: rom_data = 8'hD0;
      9'h19A: rom_data = 8'h6A;
      9'h19B: rom_data = 8'hCC;
      9'h19C: rom_data = 8'h9E;
      9'h19D: rom_data = 8'h98;
      9'h19E: rom_data = 8'h36;
      9'h19F: rom_data = 8'h71;
      9'h1A0: rom_data = 8'hA4;
      9'h1A1: rom_data = 8'hEB;
      9'h1A2: rom_data = 8'h38;
      9'h1A3: rom_data = 8'h82;
      9'h1A4: rom_data = 8'hB9;
      9'h1A5: rom_data = 8'h38;
      9'h1A6: rom_data = 8'h1F;
      9'h1A7: rom_data = 8'hC1;
      9'h1A8: rom_data = 8'hF9;
      9'h1A9: rom_data = 8'h90;
      9'h1AA: rom_data = 8'h00;
      9'h1AB: rom_data = 8'h3D;
      9'h1AC: rom_data = 8'hEB;
      9'h1AD: rom_data = 8'h10;
      9'h1AE: rom_data = 8'h76;
      9'h1AF: rom_data = 8'hAF;
      9'h1B0: rom_data = 8'h99;
      9'h1B1: rom_data = 8'hFF;
      9'h1B2: rom_data = 8'hE4;
      9'h1B3: rom_data = 8'h97;
      9'h1B4: rom_data = 8'hBF;
      9'h1B5: rom_data = 8'h57;
      9'h1B6: rom_data = 8'h0C;
      9'h1B7: rom_data = 8'h84;
      9'h1B8: rom_data = 8'hBE;
      9'h1B9: rom_data = 8'h09;
      9'h1BA: rom_data = 8'h42;
      9'h1BB: rom_data = 8'h3D;
      9'h1BC: rom_data = 8'hD5;
      9'h1BD: rom_data = 8'hC2;
      9'h1BE: rom_data = 8'h7D;
      9'h1BF: rom_data = 8'hD2;
      9'h1C0: rom_data = 8'h17;
      9'h1C1: rom_data = 8'h94;
      9'h1C2: rom_data = 8'hEA;
      9'h1C3: rom_data = 8'h88;
      9'h1C4: rom_data = 8'h31;
      9'h1C5: rom_data = 8'h55;
      9'h1C6: rom_data = 8'hFB;
      9'h1C7: rom_data = 8'hCD;
      9'h1C8: rom_data = 8'hD7;
      9'h1C9: rom_data = 8'hA3;
      9'h1CA: rom_data = 8'h05;
      9'h1CB: rom_data = 8'h94;
      9'h1CC: rom_data = 8'h99;
      9'h1CD: rom_data = 8'hB7;
      9'h1CE: rom_data = 8'h2D;
      9'h1CF: rom_data = 8'h38;
      9'h1D0: rom_data = 8'hD0;
      9'h1D1: rom_data = 8'h34;
      9'h1D2: rom_data = 8'hCE;
      9'h1D3: rom_data = 8'h2A;
      9'h1D4: rom_data = 8'hEF;
      9'h1D5: rom_data = 8'h3B;
      9'h1D6: rom_data = 8'hA0;
      9'h1D7: rom_data = 8'h3C;
      9'h1D8: rom_data = 8'h0C;
      9'h1D9: rom_data = 8'h39;
      9'h1DA: rom_data = 8'h1A;
      9'h1DB: rom_data = 8'hB4;
      9'h1DC: rom_data = 8'hFD;
      9'h1DD: rom_data = 8'hAD;
      9'h1DE: rom_data = 8'h2B;
      9'h1DF: rom_data = 8'hE6;
      9'h1E0: rom_data = 8'h70;
      9'h1E1: rom_data = 8'h7D;
      9'h1E2: rom_data = 8'h53;
      9'h1E3: rom_data = 8'h94;
      9'h1E4: rom_data = 8'h6C;
      9'h1E5: rom_data = 8'hE4;
      9'h1E6: rom_data = 8'hA5;
      9'h1E7: rom_data = 8'hC1;
      9'h1E8: rom_data = 8'h1C;
      9'h1E9: rom_data = 8'h29;
      9'h1EA: rom_data = 8'hA3;
      9'h1EB: rom_data = 8'hB1;
      9'h1EC: rom_data = 8'h28;
      9'h1ED: rom_data = 8'h51;
      9'h1EE: rom_data = 8'hDA;
      9'h1EF: rom_data = 8'h9A;
      9'h1F0: rom_data = 8'h96;
      9'h1F1: rom_data = 8'hDD;
      9'h1F2: rom_data = 8'h4B;
      9'h1F3: rom_data = 8'h7E;
      9'h1F4: rom_data = 8'h56;
      9'h1F5: rom_data = 8'hBF;
      9'h1F6: rom_data = 8'h5A;
      9'h1F7: rom_data = 8'h41;
      9'h1F8: rom_data = 8'h6B;
      9'h1F9: rom_data = 8'hFF;
      9'h1FA: rom_data = 8'h06;
      9'h1FB: rom_data = 8'hC8;
      9'h1FC: rom_data = 8'hB3;
      9'h1FD: rom_data = 8'h63;
      9'h1FE: rom_data = 8'h2E;
      9'h1FF: rom_data = 8'h17;

      default: rom_data = 8'h00;
    endcase
  end

  always @(posedge clk) begin
    if (~rst_n) begin
      rom_addr_r <= 0;
      rom_data_r <= 0;
    end else begin
      rom_addr_r <= rom_addr;
      rom_data_r <= rom_data;
    end
  end

  assign rom_addr = counter[10:2];
  assign audio_sample = {8'h00, rom_data_r};

// Audio end

  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      counter <= counter + 1;
    end
  end
  
endmodule
