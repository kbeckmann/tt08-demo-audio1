/*
 * Copyright (c) 2024 Konrad Beckmann
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_vga_example(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,   // Dedicated outputs
  input  wire [7:0] uio_in,   // IOs: Input path
  output wire [7:0] uio_out,  // IOs: Output path
  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
  input  wire       ena,      // always 1 when the design is powered, so you can ignore it
  input  wire       clk,      // clock
  input  wire       rst_n     // reset_n - low to reset
);

  // Audio signals
  wire audio_out;
  wire [15:0] audio_sample;

  // TinyVGA PMOD
  // assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};
  assign uo_out = 8'b00000000;

  // Audio PMOD
  assign uio_out = {audio_out, 7'b0000000};
  assign uio_oe = 8'b10000000;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in, uio_in};

  reg [10:0] counter;

// Audio start
  pdm #(.N(16)) pdm_gen(
    .clk(clk),
    .rst_n(rst_n),
    .pdm_in(audio_sample),
    .pdm_out(audio_out)
  );

  // ROM
  wire [9:0] rom_addr;
  reg  [9:0] rom_addr_r;
  reg  [7:0] rom_data_r;
  reg  [7:0] rom_content[1024];

  initial begin
  rom_content[0] = 8'h68;
  rom_content[1] = 8'h40;
  rom_content[2] = 8'h94;
  rom_content[3] = 8'hE0;
  rom_content[4] = 8'hF5;
  rom_content[5] = 8'h23;
  rom_content[6] = 8'h13;
  rom_content[7] = 8'h0E;
  rom_content[8] = 8'h18;
  rom_content[9] = 8'h18;
  rom_content[10] = 8'h8D;
  rom_content[11] = 8'h5A;
  rom_content[12] = 8'hB9;
  rom_content[13] = 8'hC1;
  rom_content[14] = 8'h10;
  rom_content[15] = 8'hFB;
  rom_content[16] = 8'h77;
  rom_content[17] = 8'h01;
  rom_content[18] = 8'h0D;
  rom_content[19] = 8'h19;
  rom_content[20] = 8'hA1;
  rom_content[21] = 8'hCD;
  rom_content[22] = 8'hCD;
  rom_content[23] = 8'h6B;
  rom_content[24] = 8'h3E;
  rom_content[25] = 8'h92;
  rom_content[26] = 8'hED;
  rom_content[27] = 8'h02;
  rom_content[28] = 8'h63;
  rom_content[29] = 8'hB1;
  rom_content[30] = 8'h89;
  rom_content[31] = 8'h4A;
  rom_content[32] = 8'h32;
  rom_content[33] = 8'h8F;
  rom_content[34] = 8'hF3;
  rom_content[35] = 8'h12;
  rom_content[36] = 8'h14;
  rom_content[37] = 8'hC9;
  rom_content[38] = 8'hCA;
  rom_content[39] = 8'h11;
  rom_content[40] = 8'h8F;
  rom_content[41] = 8'hE4;
  rom_content[42] = 8'h17;
  rom_content[43] = 8'h5A;
  rom_content[44] = 8'hD0;
  rom_content[45] = 8'h69;
  rom_content[46] = 8'h4D;
  rom_content[47] = 8'h09;
  rom_content[48] = 8'h05;
  rom_content[49] = 8'hF6;
  rom_content[50] = 8'h80;
  rom_content[51] = 8'h13;
  rom_content[52] = 8'h43;
  rom_content[53] = 8'hE5;
  rom_content[54] = 8'hCF;
  rom_content[55] = 8'h8E;
  rom_content[56] = 8'h91;
  rom_content[57] = 8'h1D;
  rom_content[58] = 8'hC0;
  rom_content[59] = 8'h13;
  rom_content[60] = 8'h3D;
  rom_content[61] = 8'hB1;
  rom_content[62] = 8'hB1;
  rom_content[63] = 8'h01;
  rom_content[64] = 8'h7C;
  rom_content[65] = 8'hF4;
  rom_content[66] = 8'h99;
  rom_content[67] = 8'h1E;
  rom_content[68] = 8'h1C;
  rom_content[69] = 8'h32;
  rom_content[70] = 8'h42;
  rom_content[71] = 8'h48;
  rom_content[72] = 8'hDB;
  rom_content[73] = 8'h09;
  rom_content[74] = 8'hC8;
  rom_content[75] = 8'h5D;
  rom_content[76] = 8'hF3;
  rom_content[77] = 8'hC8;
  rom_content[78] = 8'h79;
  rom_content[79] = 8'hD3;
  rom_content[80] = 8'hA7;
  rom_content[81] = 8'h92;
  rom_content[82] = 8'h66;
  rom_content[83] = 8'h39;
  rom_content[84] = 8'h92;
  rom_content[85] = 8'hC4;
  rom_content[86] = 8'h05;
  rom_content[87] = 8'hCA;
  rom_content[88] = 8'h36;
  rom_content[89] = 8'h6C;
  rom_content[90] = 8'h14;
  rom_content[91] = 8'h51;
  rom_content[92] = 8'h6E;
  rom_content[93] = 8'hA2;
  rom_content[94] = 8'hA0;
  rom_content[95] = 8'h81;
  rom_content[96] = 8'h8F;
  rom_content[97] = 8'hF0;
  rom_content[98] = 8'h60;
  rom_content[99] = 8'h7C;
  rom_content[100] = 8'h27;
  rom_content[101] = 8'h1E;
  rom_content[102] = 8'hE5;
  rom_content[103] = 8'h87;
  rom_content[104] = 8'h30;
  rom_content[105] = 8'h24;
  rom_content[106] = 8'h96;
  rom_content[107] = 8'h9F;
  rom_content[108] = 8'h65;
  rom_content[109] = 8'h34;
  rom_content[110] = 8'h96;
  rom_content[111] = 8'hF1;
  rom_content[112] = 8'h30;
  rom_content[113] = 8'hFE;
  rom_content[114] = 8'h2F;
  rom_content[115] = 8'hF1;
  rom_content[116] = 8'h1C;
  rom_content[117] = 8'hF6;
  rom_content[118] = 8'hE1;
  rom_content[119] = 8'hE1;
  rom_content[120] = 8'h75;
  rom_content[121] = 8'h7E;
  rom_content[122] = 8'hC1;
  rom_content[123] = 8'h8C;
  rom_content[124] = 8'h3E;
  rom_content[125] = 8'hB8;
  rom_content[126] = 8'h01;
  rom_content[127] = 8'h03;
  rom_content[128] = 8'h0D;
  rom_content[129] = 8'h20;
  rom_content[130] = 8'h87;
  rom_content[131] = 8'h55;
  rom_content[132] = 8'h17;
  rom_content[133] = 8'h58;
  rom_content[134] = 8'hD6;
  rom_content[135] = 8'h6A;
  rom_content[136] = 8'hD9;
  rom_content[137] = 8'hCC;
  rom_content[138] = 8'h96;
  rom_content[139] = 8'h3F;
  rom_content[140] = 8'hED;
  rom_content[141] = 8'hBF;
  rom_content[142] = 8'hB4;
  rom_content[143] = 8'hED;
  rom_content[144] = 8'h76;
  rom_content[145] = 8'hF8;
  rom_content[146] = 8'h69;
  rom_content[147] = 8'hC3;
  rom_content[148] = 8'hD6;
  rom_content[149] = 8'h1F;
  rom_content[150] = 8'hC0;
  rom_content[151] = 8'hF6;
  rom_content[152] = 8'hDF;
  rom_content[153] = 8'h92;
  rom_content[154] = 8'h0F;
  rom_content[155] = 8'h7E;
  rom_content[156] = 8'hC2;
  rom_content[157] = 8'hC5;
  rom_content[158] = 8'h8C;
  rom_content[159] = 8'hD3;
  rom_content[160] = 8'h6C;
  rom_content[161] = 8'hB2;
  rom_content[162] = 8'hC4;
  rom_content[163] = 8'h32;
  rom_content[164] = 8'h42;
  rom_content[165] = 8'hB9;
  rom_content[166] = 8'hCD;
  rom_content[167] = 8'h29;
  rom_content[168] = 8'hCF;
  rom_content[169] = 8'hCC;
  rom_content[170] = 8'hDC;
  rom_content[171] = 8'hEC;
  rom_content[172] = 8'h48;
  rom_content[173] = 8'h08;
  rom_content[174] = 8'hAA;
  rom_content[175] = 8'hA3;
  rom_content[176] = 8'h5B;
  rom_content[177] = 8'h87;
  rom_content[178] = 8'hC0;
  rom_content[179] = 8'hAA;
  rom_content[180] = 8'h98;
  rom_content[181] = 8'h5D;
  rom_content[182] = 8'h71;
  rom_content[183] = 8'h0C;
  rom_content[184] = 8'hA2;
  rom_content[185] = 8'hAC;
  rom_content[186] = 8'hB4;
  rom_content[187] = 8'hEA;
  rom_content[188] = 8'h16;
  rom_content[189] = 8'h72;
  rom_content[190] = 8'h09;
  rom_content[191] = 8'h9D;
  rom_content[192] = 8'h30;
  rom_content[193] = 8'h1A;
  rom_content[194] = 8'hE5;
  rom_content[195] = 8'hBA;
  rom_content[196] = 8'hFB;
  rom_content[197] = 8'h48;
  rom_content[198] = 8'h5B;
  rom_content[199] = 8'hD0;
  rom_content[200] = 8'hD2;
  rom_content[201] = 8'h27;
  rom_content[202] = 8'h86;
  rom_content[203] = 8'h9C;
  rom_content[204] = 8'h40;
  rom_content[205] = 8'h7B;
  rom_content[206] = 8'hAB;
  rom_content[207] = 8'h4F;
  rom_content[208] = 8'hED;
  rom_content[209] = 8'hF7;
  rom_content[210] = 8'h06;
  rom_content[211] = 8'hB5;
  rom_content[212] = 8'hF1;
  rom_content[213] = 8'h78;
  rom_content[214] = 8'h79;
  rom_content[215] = 8'hBB;
  rom_content[216] = 8'h94;
  rom_content[217] = 8'h69;
  rom_content[218] = 8'h00;
  rom_content[219] = 8'h47;
  rom_content[220] = 8'h61;
  rom_content[221] = 8'hB6;
  rom_content[222] = 8'h2A;
  rom_content[223] = 8'h6D;
  rom_content[224] = 8'hCF;
  rom_content[225] = 8'hB8;
  rom_content[226] = 8'hC6;
  rom_content[227] = 8'hDA;
  rom_content[228] = 8'h63;
  rom_content[229] = 8'h8A;
  rom_content[230] = 8'h4B;
  rom_content[231] = 8'hB8;
  rom_content[232] = 8'h13;
  rom_content[233] = 8'hDF;
  rom_content[234] = 8'h60;
  rom_content[235] = 8'hDB;
  rom_content[236] = 8'h4D;
  rom_content[237] = 8'hAF;
  rom_content[238] = 8'h9B;
  rom_content[239] = 8'h39;
  rom_content[240] = 8'hF1;
  rom_content[241] = 8'h2B;
  rom_content[242] = 8'h3D;
  rom_content[243] = 8'h32;
  rom_content[244] = 8'h0E;
  rom_content[245] = 8'hC9;
  rom_content[246] = 8'h49;
  rom_content[247] = 8'h80;
  rom_content[248] = 8'h6E;
  rom_content[249] = 8'h2A;
  rom_content[250] = 8'hE6;
  rom_content[251] = 8'h7B;
  rom_content[252] = 8'hA2;
  rom_content[253] = 8'hC4;
  rom_content[254] = 8'h42;
  rom_content[255] = 8'h91;
  rom_content[256] = 8'hA6;
  rom_content[257] = 8'hE8;
  rom_content[258] = 8'h7E;
  rom_content[259] = 8'hFB;
  rom_content[260] = 8'h3E;
  rom_content[261] = 8'hF3;
  rom_content[262] = 8'hA7;
  rom_content[263] = 8'h90;
  rom_content[264] = 8'hEB;
  rom_content[265] = 8'hFE;
  rom_content[266] = 8'hCF;
  rom_content[267] = 8'hCD;
  rom_content[268] = 8'h7D;
  rom_content[269] = 8'hAD;
  rom_content[270] = 8'h37;
  rom_content[271] = 8'h4A;
  rom_content[272] = 8'h03;
  rom_content[273] = 8'hAA;
  rom_content[274] = 8'hC3;
  rom_content[275] = 8'h92;
  rom_content[276] = 8'h6D;
  rom_content[277] = 8'h44;
  rom_content[278] = 8'h53;
  rom_content[279] = 8'h05;
  rom_content[280] = 8'h47;
  rom_content[281] = 8'h68;
  rom_content[282] = 8'h84;
  rom_content[283] = 8'h5D;
  rom_content[284] = 8'hE1;
  rom_content[285] = 8'h50;
  rom_content[286] = 8'h80;
  rom_content[287] = 8'hE9;
  rom_content[288] = 8'hB1;
  rom_content[289] = 8'h74;
  rom_content[290] = 8'hD8;
  rom_content[291] = 8'h9D;
  rom_content[292] = 8'h9E;
  rom_content[293] = 8'hEF;
  rom_content[294] = 8'h30;
  rom_content[295] = 8'h86;
  rom_content[296] = 8'h11;
  rom_content[297] = 8'h89;
  rom_content[298] = 8'h9C;
  rom_content[299] = 8'h98;
  rom_content[300] = 8'hB7;
  rom_content[301] = 8'h39;
  rom_content[302] = 8'h1D;
  rom_content[303] = 8'h7E;
  rom_content[304] = 8'hEA;
  rom_content[305] = 8'h29;
  rom_content[306] = 8'hC5;
  rom_content[307] = 8'h86;
  rom_content[308] = 8'hC0;
  rom_content[309] = 8'h75;
  rom_content[310] = 8'h9D;
  rom_content[311] = 8'hAF;
  rom_content[312] = 8'h07;
  rom_content[313] = 8'h2A;
  rom_content[314] = 8'h48;
  rom_content[315] = 8'hD4;
  rom_content[316] = 8'h35;
  rom_content[317] = 8'h48;
  rom_content[318] = 8'h00;
  rom_content[319] = 8'h3E;
  rom_content[320] = 8'h31;
  rom_content[321] = 8'hD2;
  rom_content[322] = 8'h6A;
  rom_content[323] = 8'h53;
  rom_content[324] = 8'h35;
  rom_content[325] = 8'h6C;
  rom_content[326] = 8'hE8;
  rom_content[327] = 8'h25;
  rom_content[328] = 8'h57;
  rom_content[329] = 8'h9A;
  rom_content[330] = 8'h0C;
  rom_content[331] = 8'h9C;
  rom_content[332] = 8'h99;
  rom_content[333] = 8'hA3;
  rom_content[334] = 8'h4E;
  rom_content[335] = 8'h12;
  rom_content[336] = 8'h87;
  rom_content[337] = 8'h45;
  rom_content[338] = 8'h52;
  rom_content[339] = 8'h9B;
  rom_content[340] = 8'hD0;
  rom_content[341] = 8'h16;
  rom_content[342] = 8'hF6;
  rom_content[343] = 8'hF7;
  rom_content[344] = 8'h54;
  rom_content[345] = 8'hB6;
  rom_content[346] = 8'h5A;
  rom_content[347] = 8'hF2;
  rom_content[348] = 8'h24;
  rom_content[349] = 8'h20;
  rom_content[350] = 8'h6B;
  rom_content[351] = 8'h33;
  rom_content[352] = 8'h1D;
  rom_content[353] = 8'h25;
  rom_content[354] = 8'h89;
  rom_content[355] = 8'hF5;
  rom_content[356] = 8'hAD;
  rom_content[357] = 8'hA2;
  rom_content[358] = 8'hA3;
  rom_content[359] = 8'h89;
  rom_content[360] = 8'h8D;
  rom_content[361] = 8'h2E;
  rom_content[362] = 8'h57;
  rom_content[363] = 8'hC2;
  rom_content[364] = 8'h98;
  rom_content[365] = 8'h19;
  rom_content[366] = 8'h3B;
  rom_content[367] = 8'h78;
  rom_content[368] = 8'h05;
  rom_content[369] = 8'h7B;
  rom_content[370] = 8'h70;
  rom_content[371] = 8'h37;
  rom_content[372] = 8'h59;
  rom_content[373] = 8'h4D;
  rom_content[374] = 8'h2E;
  rom_content[375] = 8'hF8;
  rom_content[376] = 8'h75;
  rom_content[377] = 8'h17;
  rom_content[378] = 8'hD3;
  rom_content[379] = 8'h8D;
  rom_content[380] = 8'h1D;
  rom_content[381] = 8'h2C;
  rom_content[382] = 8'hCE;
  rom_content[383] = 8'h9E;
  rom_content[384] = 8'hC2;
  rom_content[385] = 8'h87;
  rom_content[386] = 8'h63;
  rom_content[387] = 8'h5E;
  rom_content[388] = 8'hA7;
  rom_content[389] = 8'hB9;
  rom_content[390] = 8'h5B;
  rom_content[391] = 8'h3C;
  rom_content[392] = 8'hD9;
  rom_content[393] = 8'hCA;
  rom_content[394] = 8'hAE;
  rom_content[395] = 8'h1D;
  rom_content[396] = 8'h69;
  rom_content[397] = 8'h43;
  rom_content[398] = 8'h68;
  rom_content[399] = 8'h86;
  rom_content[400] = 8'h06;
  rom_content[401] = 8'h9C;
  rom_content[402] = 8'hB4;
  rom_content[403] = 8'h16;
  rom_content[404] = 8'h11;
  rom_content[405] = 8'h30;
  rom_content[406] = 8'h57;
  rom_content[407] = 8'h56;
  rom_content[408] = 8'h6C;
  rom_content[409] = 8'hA4;
  rom_content[410] = 8'hD8;
  rom_content[411] = 8'hAD;
  rom_content[412] = 8'hC0;
  rom_content[413] = 8'hD3;
  rom_content[414] = 8'h99;
  rom_content[415] = 8'h70;
  rom_content[416] = 8'h01;
  rom_content[417] = 8'hF9;
  rom_content[418] = 8'h57;
  rom_content[419] = 8'h9C;
  rom_content[420] = 8'hC6;
  rom_content[421] = 8'h7A;
  rom_content[422] = 8'hE7;
  rom_content[423] = 8'h60;
  rom_content[424] = 8'h8C;
  rom_content[425] = 8'hEF;
  rom_content[426] = 8'h31;
  rom_content[427] = 8'h31;
  rom_content[428] = 8'hD9;
  rom_content[429] = 8'h40;
  rom_content[430] = 8'h4B;
  rom_content[431] = 8'h79;
  rom_content[432] = 8'h09;
  rom_content[433] = 8'h3E;
  rom_content[434] = 8'hEB;
  rom_content[435] = 8'h7A;
  rom_content[436] = 8'hD3;
  rom_content[437] = 8'hAD;
  rom_content[438] = 8'h78;
  rom_content[439] = 8'h8D;
  rom_content[440] = 8'h96;
  rom_content[441] = 8'h1E;
  rom_content[442] = 8'hE1;
  rom_content[443] = 8'hDB;
  rom_content[444] = 8'hA8;
  rom_content[445] = 8'h9F;
  rom_content[446] = 8'h42;
  rom_content[447] = 8'hD6;
  rom_content[448] = 8'h19;
  rom_content[449] = 8'h18;
  rom_content[450] = 8'h83;
  rom_content[451] = 8'h99;
  rom_content[452] = 8'h82;
  rom_content[453] = 8'h9D;
  rom_content[454] = 8'hDF;
  rom_content[455] = 8'h18;
  rom_content[456] = 8'h08;
  rom_content[457] = 8'hC8;
  rom_content[458] = 8'hBC;
  rom_content[459] = 8'hE4;
  rom_content[460] = 8'h5E;
  rom_content[461] = 8'h7B;
  rom_content[462] = 8'hC5;
  rom_content[463] = 8'h34;
  rom_content[464] = 8'h25;
  rom_content[465] = 8'h6C;
  rom_content[466] = 8'h72;
  rom_content[467] = 8'h5A;
  rom_content[468] = 8'h95;
  rom_content[469] = 8'h2F;
  rom_content[470] = 8'hB2;
  rom_content[471] = 8'h78;
  rom_content[472] = 8'hC7;
  rom_content[473] = 8'h01;
  rom_content[474] = 8'h0F;
  rom_content[475] = 8'h11;
  rom_content[476] = 8'h4E;
  rom_content[477] = 8'h01;
  rom_content[478] = 8'h00;
  rom_content[479] = 8'h95;
  rom_content[480] = 8'h3C;
  rom_content[481] = 8'h6F;
  rom_content[482] = 8'h82;
  rom_content[483] = 8'h8A;
  rom_content[484] = 8'h5A;
  rom_content[485] = 8'hFB;
  rom_content[486] = 8'hD8;
  rom_content[487] = 8'hAA;
  rom_content[488] = 8'hD3;
  rom_content[489] = 8'h71;
  rom_content[490] = 8'hC9;
  rom_content[491] = 8'h59;
  rom_content[492] = 8'h89;
  rom_content[493] = 8'h8D;
  rom_content[494] = 8'h4D;
  rom_content[495] = 8'hC3;
  rom_content[496] = 8'hB6;
  rom_content[497] = 8'h6D;
  rom_content[498] = 8'hCD;
  rom_content[499] = 8'h52;
  rom_content[500] = 8'h9F;
  rom_content[501] = 8'hBF;
  rom_content[502] = 8'h43;
  rom_content[503] = 8'hF0;
  rom_content[504] = 8'hA4;
  rom_content[505] = 8'hFC;
  rom_content[506] = 8'hE0;
  rom_content[507] = 8'hB0;
  rom_content[508] = 8'h42;
  rom_content[509] = 8'h4F;
  rom_content[510] = 8'h63;
  rom_content[511] = 8'h72;
  rom_content[512] = 8'h05;
  rom_content[513] = 8'hB1;
  rom_content[514] = 8'hF2;
  rom_content[515] = 8'hB5;
  rom_content[516] = 8'hB5;
  rom_content[517] = 8'hEB;
  rom_content[518] = 8'h4D;
  rom_content[519] = 8'hB5;
  rom_content[520] = 8'h7C;
  rom_content[521] = 8'hDE;
  rom_content[522] = 8'h05;
  rom_content[523] = 8'h09;
  rom_content[524] = 8'hE4;
  rom_content[525] = 8'h04;
  rom_content[526] = 8'h80;
  rom_content[527] = 8'h73;
  rom_content[528] = 8'h05;
  rom_content[529] = 8'hE6;
  rom_content[530] = 8'hC4;
  rom_content[531] = 8'h08;
  rom_content[532] = 8'h3A;
  rom_content[533] = 8'h91;
  rom_content[534] = 8'hB4;
  rom_content[535] = 8'h3B;
  rom_content[536] = 8'hA7;
  rom_content[537] = 8'hFE;
  rom_content[538] = 8'h64;
  rom_content[539] = 8'hD2;
  rom_content[540] = 8'hFE;
  rom_content[541] = 8'h33;
  rom_content[542] = 8'h7E;
  rom_content[543] = 8'h93;
  rom_content[544] = 8'hED;
  rom_content[545] = 8'hC1;
  rom_content[546] = 8'hBE;
  rom_content[547] = 8'hC7;
  rom_content[548] = 8'h5F;
  rom_content[549] = 8'h67;
  rom_content[550] = 8'hFB;
  rom_content[551] = 8'h2D;
  rom_content[552] = 8'h7A;
  rom_content[553] = 8'hEB;
  rom_content[554] = 8'h17;
  rom_content[555] = 8'h11;
  rom_content[556] = 8'h35;
  rom_content[557] = 8'h43;
  rom_content[558] = 8'hC7;
  rom_content[559] = 8'hFD;
  rom_content[560] = 8'hC6;
  rom_content[561] = 8'hB1;
  rom_content[562] = 8'h15;
  rom_content[563] = 8'hE4;
  rom_content[564] = 8'h7C;
  rom_content[565] = 8'h4D;
  rom_content[566] = 8'h29;
  rom_content[567] = 8'h28;
  rom_content[568] = 8'h7D;
  rom_content[569] = 8'h6D;
  rom_content[570] = 8'h47;
  rom_content[571] = 8'hEC;
  rom_content[572] = 8'h7E;
  rom_content[573] = 8'h76;
  rom_content[574] = 8'hBB;
  rom_content[575] = 8'hB7;
  rom_content[576] = 8'hA1;
  rom_content[577] = 8'h2F;
  rom_content[578] = 8'h88;
  rom_content[579] = 8'hEB;
  rom_content[580] = 8'hFC;
  rom_content[581] = 8'h0E;
  rom_content[582] = 8'h7A;
  rom_content[583] = 8'h46;
  rom_content[584] = 8'h74;
  rom_content[585] = 8'hA5;
  rom_content[586] = 8'h92;
  rom_content[587] = 8'h04;
  rom_content[588] = 8'h4F;
  rom_content[589] = 8'h13;
  rom_content[590] = 8'h11;
  rom_content[591] = 8'h32;
  rom_content[592] = 8'hC5;
  rom_content[593] = 8'hD3;
  rom_content[594] = 8'h7C;
  rom_content[595] = 8'hCE;
  rom_content[596] = 8'hC3;
  rom_content[597] = 8'hB6;
  rom_content[598] = 8'h23;
  rom_content[599] = 8'hAA;
  rom_content[600] = 8'h27;
  rom_content[601] = 8'h2F;
  rom_content[602] = 8'h30;
  rom_content[603] = 8'hDE;
  rom_content[604] = 8'hD0;
  rom_content[605] = 8'h1F;
  rom_content[606] = 8'h02;
  rom_content[607] = 8'h8D;
  rom_content[608] = 8'h10;
  rom_content[609] = 8'hB7;
  rom_content[610] = 8'h87;
  rom_content[611] = 8'h1B;
  rom_content[612] = 8'hCF;
  rom_content[613] = 8'h9A;
  rom_content[614] = 8'h9A;
  rom_content[615] = 8'h99;
  rom_content[616] = 8'h88;
  rom_content[617] = 8'hAC;
  rom_content[618] = 8'h6A;
  rom_content[619] = 8'h1B;
  rom_content[620] = 8'h7C;
  rom_content[621] = 8'hA9;
  rom_content[622] = 8'hB2;
  rom_content[623] = 8'h96;
  rom_content[624] = 8'h9F;
  rom_content[625] = 8'hF8;
  rom_content[626] = 8'h75;
  rom_content[627] = 8'h8D;
  rom_content[628] = 8'hB8;
  rom_content[629] = 8'h56;
  rom_content[630] = 8'h80;
  rom_content[631] = 8'h9E;
  rom_content[632] = 8'h9E;
  rom_content[633] = 8'h10;
  rom_content[634] = 8'h78;
  rom_content[635] = 8'h74;
  rom_content[636] = 8'hE1;
  rom_content[637] = 8'h5B;
  rom_content[638] = 8'h66;
  rom_content[639] = 8'hB8;
  rom_content[640] = 8'hDB;
  rom_content[641] = 8'hAA;
  rom_content[642] = 8'h1A;
  rom_content[643] = 8'h0E;
  rom_content[644] = 8'hC9;
  rom_content[645] = 8'hDA;
  rom_content[646] = 8'hE1;
  rom_content[647] = 8'hE4;
  rom_content[648] = 8'h24;
  rom_content[649] = 8'hEF;
  rom_content[650] = 8'hCF;
  rom_content[651] = 8'hD9;
  rom_content[652] = 8'h98;
  rom_content[653] = 8'hB2;
  rom_content[654] = 8'h30;
  rom_content[655] = 8'h64;
  rom_content[656] = 8'h0E;
  rom_content[657] = 8'h1C;
  rom_content[658] = 8'hFB;
  rom_content[659] = 8'h33;
  rom_content[660] = 8'h25;
  rom_content[661] = 8'hDE;
  rom_content[662] = 8'h67;
  rom_content[663] = 8'h19;
  rom_content[664] = 8'h63;
  rom_content[665] = 8'hD8;
  rom_content[666] = 8'hC3;
  rom_content[667] = 8'h9A;
  rom_content[668] = 8'h0E;
  rom_content[669] = 8'h88;
  rom_content[670] = 8'hB3;
  rom_content[671] = 8'hA0;
  rom_content[672] = 8'h44;
  rom_content[673] = 8'hFD;
  rom_content[674] = 8'hB3;
  rom_content[675] = 8'h3C;
  rom_content[676] = 8'h43;
  rom_content[677] = 8'h34;
  rom_content[678] = 8'h5A;
  rom_content[679] = 8'hBC;
  rom_content[680] = 8'h46;
  rom_content[681] = 8'h7F;
  rom_content[682] = 8'h9B;
  rom_content[683] = 8'hF1;
  rom_content[684] = 8'h58;
  rom_content[685] = 8'hC9;
  rom_content[686] = 8'h92;
  rom_content[687] = 8'h69;
  rom_content[688] = 8'h4A;
  rom_content[689] = 8'h36;
  rom_content[690] = 8'h05;
  rom_content[691] = 8'hD2;
  rom_content[692] = 8'h36;
  rom_content[693] = 8'hA6;
  rom_content[694] = 8'hB6;
  rom_content[695] = 8'h0A;
  rom_content[696] = 8'h07;
  rom_content[697] = 8'h96;
  rom_content[698] = 8'h6D;
  rom_content[699] = 8'hE4;
  rom_content[700] = 8'h9F;
  rom_content[701] = 8'h95;
  rom_content[702] = 8'hBF;
  rom_content[703] = 8'hB3;
  rom_content[704] = 8'hF6;
  rom_content[705] = 8'h06;
  rom_content[706] = 8'hEA;
  rom_content[707] = 8'h03;
  rom_content[708] = 8'h91;
  rom_content[709] = 8'h68;
  rom_content[710] = 8'hB0;
  rom_content[711] = 8'h3B;
  rom_content[712] = 8'h87;
  rom_content[713] = 8'h0A;
  rom_content[714] = 8'h31;
  rom_content[715] = 8'h1F;
  rom_content[716] = 8'hB4;
  rom_content[717] = 8'hEA;
  rom_content[718] = 8'hED;
  rom_content[719] = 8'h1C;
  rom_content[720] = 8'hA7;
  rom_content[721] = 8'h42;
  rom_content[722] = 8'hCB;
  rom_content[723] = 8'hB8;
  rom_content[724] = 8'hBA;
  rom_content[725] = 8'hA7;
  rom_content[726] = 8'h7A;
  rom_content[727] = 8'hDA;
  rom_content[728] = 8'h32;
  rom_content[729] = 8'h92;
  rom_content[730] = 8'hEC;
  rom_content[731] = 8'h23;
  rom_content[732] = 8'h0D;
  rom_content[733] = 8'h69;
  rom_content[734] = 8'h1E;
  rom_content[735] = 8'h00;
  rom_content[736] = 8'hF3;
  rom_content[737] = 8'h47;
  rom_content[738] = 8'hC3;
  rom_content[739] = 8'hFC;
  rom_content[740] = 8'h06;
  rom_content[741] = 8'h3F;
  rom_content[742] = 8'h98;
  rom_content[743] = 8'hB9;
  rom_content[744] = 8'h36;
  rom_content[745] = 8'h5E;
  rom_content[746] = 8'h12;
  rom_content[747] = 8'hC9;
  rom_content[748] = 8'hF7;
  rom_content[749] = 8'h5C;
  rom_content[750] = 8'hA2;
  rom_content[751] = 8'hA0;
  rom_content[752] = 8'h73;
  rom_content[753] = 8'h19;
  rom_content[754] = 8'h1C;
  rom_content[755] = 8'h28;
  rom_content[756] = 8'h0C;
  rom_content[757] = 8'hB5;
  rom_content[758] = 8'hD2;
  rom_content[759] = 8'h8A;
  rom_content[760] = 8'hF3;
  rom_content[761] = 8'h72;
  rom_content[762] = 8'h03;
  rom_content[763] = 8'h55;
  rom_content[764] = 8'hF6;
  rom_content[765] = 8'h5B;
  rom_content[766] = 8'hE3;
  rom_content[767] = 8'h6C;
  rom_content[768] = 8'h5E;
  rom_content[769] = 8'h97;
  rom_content[770] = 8'h0A;
  rom_content[771] = 8'hF6;
  rom_content[772] = 8'h6F;
  rom_content[773] = 8'hE8;
  rom_content[774] = 8'hC6;
  rom_content[775] = 8'hAA;
  rom_content[776] = 8'hC7;
  rom_content[777] = 8'h20;
  rom_content[778] = 8'h9A;
  rom_content[779] = 8'hE3;
  rom_content[780] = 8'h6C;
  rom_content[781] = 8'h3B;
  rom_content[782] = 8'hF5;
  rom_content[783] = 8'h5D;
  rom_content[784] = 8'h10;
  rom_content[785] = 8'hD3;
  rom_content[786] = 8'hBF;
  rom_content[787] = 8'h60;
  rom_content[788] = 8'hC8;
  rom_content[789] = 8'h9A;
  rom_content[790] = 8'h8B;
  rom_content[791] = 8'hAC;
  rom_content[792] = 8'h03;
  rom_content[793] = 8'hFD;
  rom_content[794] = 8'h23;
  rom_content[795] = 8'h2F;
  rom_content[796] = 8'hAE;
  rom_content[797] = 8'h79;
  rom_content[798] = 8'hDC;
  rom_content[799] = 8'h35;
  rom_content[800] = 8'hB9;
  rom_content[801] = 8'h0A;
  rom_content[802] = 8'h96;
  rom_content[803] = 8'hA6;
  rom_content[804] = 8'hC7;
  rom_content[805] = 8'hAE;
  rom_content[806] = 8'hDB;
  rom_content[807] = 8'h72;
  rom_content[808] = 8'hE6;
  rom_content[809] = 8'hF9;
  rom_content[810] = 8'hE9;
  rom_content[811] = 8'hF8;
  rom_content[812] = 8'h9E;
  rom_content[813] = 8'hD8;
  rom_content[814] = 8'h36;
  rom_content[815] = 8'h58;
  rom_content[816] = 8'h1E;
  rom_content[817] = 8'h00;
  rom_content[818] = 8'h3A;
  rom_content[819] = 8'hA3;
  rom_content[820] = 8'h4D;
  rom_content[821] = 8'h48;
  rom_content[822] = 8'hA1;
  rom_content[823] = 8'h38;
  rom_content[824] = 8'hEF;
  rom_content[825] = 8'h7C;
  rom_content[826] = 8'h39;
  rom_content[827] = 8'h35;
  rom_content[828] = 8'h68;
  rom_content[829] = 8'h75;
  rom_content[830] = 8'h8A;
  rom_content[831] = 8'hAD;
  rom_content[832] = 8'h4E;
  rom_content[833] = 8'hC6;
  rom_content[834] = 8'h19;
  rom_content[835] = 8'hEA;
  rom_content[836] = 8'h6A;
  rom_content[837] = 8'h6D;
  rom_content[838] = 8'h96;
  rom_content[839] = 8'h73;
  rom_content[840] = 8'hFC;
  rom_content[841] = 8'h6F;
  rom_content[842] = 8'h4F;
  rom_content[843] = 8'h7D;
  rom_content[844] = 8'hB7;
  rom_content[845] = 8'h21;
  rom_content[846] = 8'h23;
  rom_content[847] = 8'hE3;
  rom_content[848] = 8'hB0;
  rom_content[849] = 8'h75;
  rom_content[850] = 8'h2B;
  rom_content[851] = 8'hC4;
  rom_content[852] = 8'h14;
  rom_content[853] = 8'h9F;
  rom_content[854] = 8'h11;
  rom_content[855] = 8'h5D;
  rom_content[856] = 8'hDC;
  rom_content[857] = 8'h9E;
  rom_content[858] = 8'h91;
  rom_content[859] = 8'h0A;
  rom_content[860] = 8'hD3;
  rom_content[861] = 8'h32;
  rom_content[862] = 8'h72;
  rom_content[863] = 8'h26;
  rom_content[864] = 8'hE4;
  rom_content[865] = 8'h08;
  rom_content[866] = 8'h90;
  rom_content[867] = 8'hC0;
  rom_content[868] = 8'hA4;
  rom_content[869] = 8'h4B;
  rom_content[870] = 8'h3D;
  rom_content[871] = 8'hA4;
  rom_content[872] = 8'h4D;
  rom_content[873] = 8'h7F;
  rom_content[874] = 8'hE4;
  rom_content[875] = 8'h9F;
  rom_content[876] = 8'hEA;
  rom_content[877] = 8'h1E;
  rom_content[878] = 8'hC3;
  rom_content[879] = 8'h98;
  rom_content[880] = 8'h55;
  rom_content[881] = 8'h31;
  rom_content[882] = 8'h66;
  rom_content[883] = 8'hA5;
  rom_content[884] = 8'hEF;
  rom_content[885] = 8'hFB;
  rom_content[886] = 8'hCC;
  rom_content[887] = 8'h92;
  rom_content[888] = 8'h7F;
  rom_content[889] = 8'h19;
  rom_content[890] = 8'h72;
  rom_content[891] = 8'hCC;
  rom_content[892] = 8'h10;
  rom_content[893] = 8'h87;
  rom_content[894] = 8'h07;
  rom_content[895] = 8'h02;
  rom_content[896] = 8'hF6;
  rom_content[897] = 8'hAB;
  rom_content[898] = 8'hAC;
  rom_content[899] = 8'h02;
  rom_content[900] = 8'hA6;
  rom_content[901] = 8'hAA;
  rom_content[902] = 8'hD8;
  rom_content[903] = 8'hC4;
  rom_content[904] = 8'h0B;
  rom_content[905] = 8'hE6;
  rom_content[906] = 8'h1E;
  rom_content[907] = 8'hDE;
  rom_content[908] = 8'h4C;
  rom_content[909] = 8'hCC;
  rom_content[910] = 8'hD0;
  rom_content[911] = 8'hFC;
  rom_content[912] = 8'h8B;
  rom_content[913] = 8'hDD;
  rom_content[914] = 8'h7E;
  rom_content[915] = 8'hFB;
  rom_content[916] = 8'hF5;
  rom_content[917] = 8'h20;
  rom_content[918] = 8'hDE;
  rom_content[919] = 8'h9C;
  rom_content[920] = 8'hE1;
  rom_content[921] = 8'h98;
  rom_content[922] = 8'hF6;
  rom_content[923] = 8'hFE;
  rom_content[924] = 8'h81;
  rom_content[925] = 8'hAB;
  rom_content[926] = 8'hAE;
  rom_content[927] = 8'h38;
  rom_content[928] = 8'hDE;
  rom_content[929] = 8'h46;
  rom_content[930] = 8'hB6;
  rom_content[931] = 8'h3F;
  rom_content[932] = 8'h63;
  rom_content[933] = 8'h47;
  rom_content[934] = 8'hEF;
  rom_content[935] = 8'hF8;
  rom_content[936] = 8'h16;
  rom_content[937] = 8'h4C;
  rom_content[938] = 8'hFB;
  rom_content[939] = 8'hC6;
  rom_content[940] = 8'h4B;
  rom_content[941] = 8'h9B;
  rom_content[942] = 8'h0D;
  rom_content[943] = 8'h70;
  rom_content[944] = 8'h7D;
  rom_content[945] = 8'h81;
  rom_content[946] = 8'h6D;
  rom_content[947] = 8'h24;
  rom_content[948] = 8'h3A;
  rom_content[949] = 8'h61;
  rom_content[950] = 8'hD2;
  rom_content[951] = 8'h92;
  rom_content[952] = 8'h5B;
  rom_content[953] = 8'hB9;
  rom_content[954] = 8'h9B;
  rom_content[955] = 8'hE2;
  rom_content[956] = 8'h07;
  rom_content[957] = 8'h94;
  rom_content[958] = 8'h27;
  rom_content[959] = 8'hD2;
  rom_content[960] = 8'hBC;
  rom_content[961] = 8'hC3;
  rom_content[962] = 8'hAF;
  rom_content[963] = 8'h7C;
  rom_content[964] = 8'h07;
  rom_content[965] = 8'h8D;
  rom_content[966] = 8'hD2;
  rom_content[967] = 8'h24;
  rom_content[968] = 8'h9A;
  rom_content[969] = 8'hB7;
  rom_content[970] = 8'hA4;
  rom_content[971] = 8'h46;
  rom_content[972] = 8'hAC;
  rom_content[973] = 8'hBF;
  rom_content[974] = 8'h48;
  rom_content[975] = 8'h07;
  rom_content[976] = 8'hD9;
  rom_content[977] = 8'hAD;
  rom_content[978] = 8'hDB;
  rom_content[979] = 8'h04;
  rom_content[980] = 8'hBD;
  rom_content[981] = 8'h06;
  rom_content[982] = 8'hD9;
  rom_content[983] = 8'hE2;
  rom_content[984] = 8'h90;
  rom_content[985] = 8'hF0;
  rom_content[986] = 8'hAC;
  rom_content[987] = 8'h97;
  rom_content[988] = 8'hDA;
  rom_content[989] = 8'hE3;
  rom_content[990] = 8'h58;
  rom_content[991] = 8'h58;
  rom_content[992] = 8'h13;
  rom_content[993] = 8'h02;
  rom_content[994] = 8'hD9;
  rom_content[995] = 8'hE2;
  rom_content[996] = 8'hCD;
  rom_content[997] = 8'h7A;
  rom_content[998] = 8'h22;
  rom_content[999] = 8'hD8;
  rom_content[1000] = 8'hB6;
  rom_content[1001] = 8'hCF;
  rom_content[1002] = 8'h5F;
  rom_content[1003] = 8'h9F;
  rom_content[1004] = 8'h01;
  rom_content[1005] = 8'h40;
  rom_content[1006] = 8'h62;
  rom_content[1007] = 8'h69;
  rom_content[1008] = 8'h58;
  rom_content[1009] = 8'hCA;
  rom_content[1010] = 8'h46;
  rom_content[1011] = 8'h66;
  rom_content[1012] = 8'h4E;
  rom_content[1013] = 8'h1B;
  rom_content[1014] = 8'hDA;
  rom_content[1015] = 8'h17;
  rom_content[1016] = 8'hD9;
  rom_content[1017] = 8'hFB;
  rom_content[1018] = 8'hD9;
  rom_content[1019] = 8'hA1;
  rom_content[1020] = 8'hF6;
  rom_content[1021] = 8'h09;
  rom_content[1022] = 8'hD4;
  rom_content[1023] = 8'h8F;

  end

  always @(posedge clk) begin
    if (~rst_n) begin
      rom_addr_r <= 0;
      rom_data_r <= 0;
    end else begin
      rom_addr_r <= rom_addr;
      rom_data_r <= rom_content[rom_addr_r];
    end
  end

  assign rom_addr = counter[10:1];
  assign audio_sample = {8'h00, rom_data_r};

// Audio end

  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      counter <= counter + 1;
    end
  end
  
endmodule
